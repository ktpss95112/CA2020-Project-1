`ifndef HAZARD_DETECTION_V
`define HAZARD_DETECTION_V

module Hazard_Detection (
    Stall_o
);

output  Stall_o;

endmodule

`endif
